--------------------------------------------------------------------------------
-- Company: 
-- Engineer: Aastha Dave
--
-- Create Date:   15:42:59 05/08/2023
-- Design Name:   
-- Module Name:   /home/ise/vhdl/submit/direct/tb_addop.vhd
-- Project Name:  idea
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: addop
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb_addop IS
END tb_addop;
 
ARCHITECTURE behavior OF tb_addop IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT addop
    PORT(
         a : IN  std_logic_vector(15 downto 0);
         b : IN  std_logic_vector(15 downto 0);
         sum : OUT  std_logic_vector(15 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal a : std_logic_vector(15 downto 0) := (others => '0');
   signal b : std_logic_vector(15 downto 0) := (others => '0');

 	--Outputs
   signal sum : std_logic_vector(15 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: addop PORT MAP (
          a => a,
          b => b,
          sum => sum
        );

   -- Stimulus process
   stim_proc: process
   begin		
		a <= x"0000";
		b <= x"0000";
		wait for 10 ns;
		
		a <= x"7ce3";
		b <= x"0000";
		wait for 10 ns;
		
		a <= x"7ce3";
		b <= x"2db6";
		wait for 10 ns;

		a <= x"fce3";
		b <= x"2db6";
		wait for 10 ns;
		
		a <= x"fce3";
		b <= x"edb6";
		wait for 10 ns;
		
		a <= x"7ce3";
		b <= x"edb6";
      wait;
   end process;

END;
